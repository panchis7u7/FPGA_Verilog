module Top (x1, x2, x3, z1, z2);
input x1, x2, x3;
output z1, z2;

endmodule